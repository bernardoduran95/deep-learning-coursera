--MEF Transmisor UART: 11 Estados: Idle (1) Start (0) D0-D7 (Datos) End(0)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mef_tx_uart is

	port (

		clk	: in std_logic;	--Reloj de entrada (9600 baudios)
		rst	: in std_logic;	--Reset
		dato	: in std_logic_vector (7 downto 0) := x"00";	--Dato que se envía (8 bits, cambia 11 veces mas lento que el clock)
		tx		: out std_logic	--Señal de tx

	);

end mef_tx_uart;

architecture arch_mef_tx_uart of mef_tx_uart is

	type mef is (idle, start, d0, d1, d2, d3, d4, d5, d6, d7, stop);
	signal estado : mef;

begin

	process (clk, rst) --Con cada flanco ascendente de reloj cambio de estado
	begin

			if rst = '1' then
				
				estado <= idle;

			elsif rising_edge (clk) then

				case estado is

					when idle => estado <= start;
					when start => estado <= d0;
					when d0 => estado <= d1;
					when d1 => estado <= d2;
					when d2 => estado <= d3;
					when d3 => estado <= d4;
					when d4 => estado <= d5;
					when d5 => estado <= d6;
					when d6 => estado <= d7;
					when d7 => estado <= stop;
					when stop => estado <= idle;

				end case;

			end if;

	end process;
	
	process (estado, dato) --Cada vez que cambia el estado o el dato envío el bit correspondiente
	begin

			case estado is

				when idle => tx <= '1';
				when start => tx <= '0';
				when d0 => tx <= dato(0);
				when d1 => tx <= dato(1);
				when d2 => tx <= dato(2);
				when d3 => tx <= dato(3);
				when d4 => tx <= dato(4);
				when d5 => tx <= dato(5);
				when d6 => tx <= dato(6);
				when d7 => tx <= dato(7);
				when stop => tx <= '0';

			end case;

	end process;

end arch_mef_tx_uart;